// mse.v

// Generated using ACDS version 12.1sp1 243 at 2013.07.21.16:14:45

`timescale 1 ps / 1 ps
module mse (
		output wire  qsys_serial_host_0_sdo,   // qsys_serial_host_0.sdo
		input  wire  qsys_serial_host_0_sdi,   //                   .sdi
		input  wire  qsys_serial_host_0_clk,   //                   .clk
		input  wire  qsys_serial_host_0_sle,   //                   .sle
		output wire  qsys_serial_host_0_srdy,  //                   .srdy
		input  wire  qsys_serial_host_0_reset  //                   .reset
	);

	wire         qsys_serial_host_0_mrst_reset;                                                            // qsys_serial_host_0:rso_MRST_reset -> [addr_router:reset, basic_SysID_0:rsi_MRST_reset, basic_SysID_0_SysID_translator:reset, basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:reset, basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux:reset, id_router:reset, id_router_001:reset, limiter:reset, qsys_serial_host_0_m1_translator:reset, qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_mux:reset, test_RegRW32_0:rsi_MRST_reset, test_RegRW32_0_test_translator:reset, test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:reset, test_RegRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         qsys_serial_host_0_mclk_clk;                                                              // qsys_serial_host_0:cso_MCLK_clk -> [addr_router:clk, basic_SysID_0:csi_MCLK_clk, basic_SysID_0_SysID_translator:clk, basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:clk, basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cmd_xbar_demux:clk, id_router:clk, id_router_001:clk, limiter:clk, qsys_serial_host_0_m1_translator:clk, qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_mux:clk, test_RegRW32_0:csi_MCLK_clk, test_RegRW32_0_test_translator:clk, test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:clk, test_RegRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:clk]
	wire         qsys_serial_host_0_m1_waitrequest;                                                        // qsys_serial_host_0_m1_translator:av_waitrequest -> qsys_serial_host_0:avm_M1_waitrequest
	wire   [7:0] qsys_serial_host_0_m1_address;                                                            // qsys_serial_host_0:avm_M1_address -> qsys_serial_host_0_m1_translator:av_address
	wire  [31:0] qsys_serial_host_0_m1_writedata;                                                          // qsys_serial_host_0:avm_M1_writedata -> qsys_serial_host_0_m1_translator:av_writedata
	wire         qsys_serial_host_0_m1_write;                                                              // qsys_serial_host_0:avm_M1_write -> qsys_serial_host_0_m1_translator:av_write
	wire         qsys_serial_host_0_m1_read;                                                               // qsys_serial_host_0:avm_M1_read -> qsys_serial_host_0_m1_translator:av_read
	wire  [31:0] qsys_serial_host_0_m1_readdata;                                                           // qsys_serial_host_0_m1_translator:av_readdata -> qsys_serial_host_0:avm_M1_readdata
	wire         qsys_serial_host_0_m1_begintransfer;                                                      // qsys_serial_host_0:avm_M1_begintransfer -> qsys_serial_host_0_m1_translator:av_begintransfer
	wire         qsys_serial_host_0_m1_readdatavalid;                                                      // qsys_serial_host_0_m1_translator:av_readdatavalid -> qsys_serial_host_0:avm_M1_readdatavalid
	wire   [3:0] qsys_serial_host_0_m1_byteenable;                                                         // qsys_serial_host_0:avm_M1_byteenable -> qsys_serial_host_0_m1_translator:av_byteenable
	wire         basic_sysid_0_sysid_translator_avalon_anti_slave_0_waitrequest;                           // basic_SysID_0:avs_SysID_waitrequest -> basic_SysID_0_SysID_translator:av_waitrequest
	wire   [1:0] basic_sysid_0_sysid_translator_avalon_anti_slave_0_address;                               // basic_SysID_0_SysID_translator:av_address -> basic_SysID_0:avs_SysID_address
	wire         basic_sysid_0_sysid_translator_avalon_anti_slave_0_read;                                  // basic_SysID_0_SysID_translator:av_read -> basic_SysID_0:avs_SysID_read
	wire  [31:0] basic_sysid_0_sysid_translator_avalon_anti_slave_0_readdata;                              // basic_SysID_0:avs_SysID_readdata -> basic_SysID_0_SysID_translator:av_readdata
	wire         test_regrw32_0_test_translator_avalon_anti_slave_0_waitrequest;                           // test_RegRW32_0:avs_test_waitrequest -> test_RegRW32_0_test_translator:av_waitrequest
	wire  [31:0] test_regrw32_0_test_translator_avalon_anti_slave_0_writedata;                             // test_RegRW32_0_test_translator:av_writedata -> test_RegRW32_0:avs_test_writedata
	wire         test_regrw32_0_test_translator_avalon_anti_slave_0_write;                                 // test_RegRW32_0_test_translator:av_write -> test_RegRW32_0:avs_test_write
	wire         test_regrw32_0_test_translator_avalon_anti_slave_0_read;                                  // test_RegRW32_0_test_translator:av_read -> test_RegRW32_0:avs_test_read
	wire  [31:0] test_regrw32_0_test_translator_avalon_anti_slave_0_readdata;                              // test_RegRW32_0:avs_test_readdata -> test_RegRW32_0_test_translator:av_readdata
	wire   [3:0] test_regrw32_0_test_translator_avalon_anti_slave_0_byteenable;                            // test_RegRW32_0_test_translator:av_byteenable -> test_RegRW32_0:avs_test_byteenable
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_waitrequest;                   // qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:av_waitrequest -> qsys_serial_host_0_m1_translator:uav_waitrequest
	wire   [2:0] qsys_serial_host_0_m1_translator_avalon_universal_master_0_burstcount;                    // qsys_serial_host_0_m1_translator:uav_burstcount -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] qsys_serial_host_0_m1_translator_avalon_universal_master_0_writedata;                     // qsys_serial_host_0_m1_translator:uav_writedata -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:av_writedata
	wire   [9:0] qsys_serial_host_0_m1_translator_avalon_universal_master_0_address;                       // qsys_serial_host_0_m1_translator:uav_address -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:av_address
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_lock;                          // qsys_serial_host_0_m1_translator:uav_lock -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:av_lock
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_write;                         // qsys_serial_host_0_m1_translator:uav_write -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:av_write
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_read;                          // qsys_serial_host_0_m1_translator:uav_read -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] qsys_serial_host_0_m1_translator_avalon_universal_master_0_readdata;                      // qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:av_readdata -> qsys_serial_host_0_m1_translator:uav_readdata
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_debugaccess;                   // qsys_serial_host_0_m1_translator:uav_debugaccess -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] qsys_serial_host_0_m1_translator_avalon_universal_master_0_byteenable;                    // qsys_serial_host_0_m1_translator:uav_byteenable -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:av_byteenable
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_readdatavalid;                 // qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:av_readdatavalid -> qsys_serial_host_0_m1_translator:uav_readdatavalid
	wire         basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // basic_SysID_0_SysID_translator:uav_waitrequest -> basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_burstcount;              // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:m0_burstcount -> basic_SysID_0_SysID_translator:uav_burstcount
	wire  [31:0] basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_writedata;               // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:m0_writedata -> basic_SysID_0_SysID_translator:uav_writedata
	wire   [9:0] basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_address;                 // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:m0_address -> basic_SysID_0_SysID_translator:uav_address
	wire         basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_write;                   // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:m0_write -> basic_SysID_0_SysID_translator:uav_write
	wire         basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_lock;                    // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:m0_lock -> basic_SysID_0_SysID_translator:uav_lock
	wire         basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_read;                    // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:m0_read -> basic_SysID_0_SysID_translator:uav_read
	wire  [31:0] basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_readdata;                // basic_SysID_0_SysID_translator:uav_readdata -> basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // basic_SysID_0_SysID_translator:uav_readdatavalid -> basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:m0_debugaccess -> basic_SysID_0_SysID_translator:uav_debugaccess
	wire   [3:0] basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_byteenable;              // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:m0_byteenable -> basic_SysID_0_SysID_translator:uav_byteenable
	wire         basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rf_source_valid;            // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:rf_source_valid -> basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [79:0] basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rf_source_data;             // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:rf_source_data -> basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rf_source_ready;            // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [79:0] basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:rf_sink_ready -> basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // test_RegRW32_0_test_translator:uav_waitrequest -> test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_burstcount;              // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:m0_burstcount -> test_RegRW32_0_test_translator:uav_burstcount
	wire  [31:0] test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_writedata;               // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:m0_writedata -> test_RegRW32_0_test_translator:uav_writedata
	wire   [9:0] test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_address;                 // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:m0_address -> test_RegRW32_0_test_translator:uav_address
	wire         test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_write;                   // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:m0_write -> test_RegRW32_0_test_translator:uav_write
	wire         test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_lock;                    // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:m0_lock -> test_RegRW32_0_test_translator:uav_lock
	wire         test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_read;                    // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:m0_read -> test_RegRW32_0_test_translator:uav_read
	wire  [31:0] test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_readdata;                // test_RegRW32_0_test_translator:uav_readdata -> test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // test_RegRW32_0_test_translator:uav_readdatavalid -> test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:m0_debugaccess -> test_RegRW32_0_test_translator:uav_debugaccess
	wire   [3:0] test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_byteenable;              // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:m0_byteenable -> test_RegRW32_0_test_translator:uav_byteenable
	wire         test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> test_RegRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_valid;            // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:rf_source_valid -> test_RegRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> test_RegRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [79:0] test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_data;             // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:rf_source_data -> test_RegRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_ready;            // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [79:0] test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:rf_sink_ready -> test_RegRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_endofpacket;          // qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_valid;                // qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_startofpacket;        // qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [78:0] qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_data;                 // qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_ready;                // addr_router:sink_ready -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:cp_ready
	wire         basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rp_valid;                   // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [78:0] basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rp_data;                    // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router:sink_ready -> basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:rp_ready
	wire         test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rp_valid;                   // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [78:0] test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rp_data;                    // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_001:sink_ready -> test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_src_endofpacket;                                                              // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_src_valid;                                                                    // addr_router:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_src_startofpacket;                                                            // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [78:0] addr_router_src_data;                                                                     // addr_router:src_data -> limiter:cmd_sink_data
	wire   [1:0] addr_router_src_channel;                                                                  // addr_router:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_src_ready;                                                                    // limiter:cmd_sink_ready -> addr_router:src_ready
	wire         limiter_rsp_src_endofpacket;                                                              // limiter:rsp_src_endofpacket -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                    // limiter:rsp_src_valid -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                            // limiter:rsp_src_startofpacket -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [78:0] limiter_rsp_src_data;                                                                     // limiter:rsp_src_data -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:rp_data
	wire   [1:0] limiter_rsp_src_channel;                                                                  // limiter:rsp_src_channel -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                    // qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         cmd_xbar_demux_src0_endofpacket;                                                          // cmd_xbar_demux:src0_endofpacket -> basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                // cmd_xbar_demux:src0_valid -> basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                        // cmd_xbar_demux:src0_startofpacket -> basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [78:0] cmd_xbar_demux_src0_data;                                                                 // cmd_xbar_demux:src0_data -> basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:cp_data
	wire   [1:0] cmd_xbar_demux_src0_channel;                                                              // cmd_xbar_demux:src0_channel -> basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src1_endofpacket;                                                          // cmd_xbar_demux:src1_endofpacket -> test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                // cmd_xbar_demux:src1_valid -> test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                        // cmd_xbar_demux:src1_startofpacket -> test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [78:0] cmd_xbar_demux_src1_data;                                                                 // cmd_xbar_demux:src1_data -> test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:cp_data
	wire   [1:0] cmd_xbar_demux_src1_channel;                                                              // cmd_xbar_demux:src1_channel -> test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                          // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                        // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [78:0] rsp_xbar_demux_src0_data;                                                                 // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [1:0] rsp_xbar_demux_src0_channel;                                                              // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                      // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                            // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                    // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [78:0] rsp_xbar_demux_001_src0_data;                                                             // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [1:0] rsp_xbar_demux_001_src0_channel;                                                          // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                            // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         limiter_cmd_src_endofpacket;                                                              // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                            // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [78:0] limiter_cmd_src_data;                                                                     // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [1:0] limiter_cmd_src_channel;                                                                  // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire         limiter_cmd_src_ready;                                                                    // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                             // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                   // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                           // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [78:0] rsp_xbar_mux_src_data;                                                                    // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [1:0] rsp_xbar_mux_src_channel;                                                                 // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_src_ready;                                                                   // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire         cmd_xbar_demux_src0_ready;                                                                // basic_SysID_0_SysID_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src0_ready
	wire         id_router_src_endofpacket;                                                                // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                      // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                              // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [78:0] id_router_src_data;                                                                       // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [1:0] id_router_src_channel;                                                                    // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                      // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_demux_src1_ready;                                                                // test_RegRW32_0_test_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src1_ready
	wire         id_router_001_src_endofpacket;                                                            // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                  // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                          // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [78:0] id_router_001_src_data;                                                                   // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [1:0] id_router_001_src_channel;                                                                // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                  // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire   [1:0] limiter_cmd_valid_data;                                                                   // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid

	qsys_serial_host #(
		.initial_state (9'b000000000)
	) qsys_serial_host_0 (
		.rso_MRST_reset       (qsys_serial_host_0_mrst_reset),       //        mrst.reset
		.cso_MCLK_clk         (qsys_serial_host_0_mclk_clk),         //        mclk.clk
		.avm_M1_writedata     (qsys_serial_host_0_m1_writedata),     //          m1.writedata
		.avm_M1_readdata      (qsys_serial_host_0_m1_readdata),      //            .readdata
		.avm_M1_address       (qsys_serial_host_0_m1_address),       //            .address
		.avm_M1_byteenable    (qsys_serial_host_0_m1_byteenable),    //            .byteenable
		.avm_M1_write         (qsys_serial_host_0_m1_write),         //            .write
		.avm_M1_read          (qsys_serial_host_0_m1_read),          //            .read
		.avm_M1_begintransfer (qsys_serial_host_0_m1_begintransfer), //            .begintransfer
		.avm_M1_readdatavalid (qsys_serial_host_0_m1_readdatavalid), //            .readdatavalid
		.avm_M1_waitrequest   (qsys_serial_host_0_m1_waitrequest),   //            .waitrequest
		.sdo                  (qsys_serial_host_0_sdo),              // conduit_end.export
		.sdi                  (qsys_serial_host_0_sdi),              //            .export
		.clk                  (qsys_serial_host_0_clk),              //            .export
		.sle                  (qsys_serial_host_0_sle),              //            .export
		.srdy                 (qsys_serial_host_0_srdy),             //            .export
		.reset                (qsys_serial_host_0_reset)             //            .export
	);

	basic_SysID basic_sysid_0 (
		.rsi_MRST_reset        (qsys_serial_host_0_mrst_reset),                                  //  MRST.reset
		.csi_MCLK_clk          (qsys_serial_host_0_mclk_clk),                                    //  MCLK.clk
		.avs_SysID_readdata    (basic_sysid_0_sysid_translator_avalon_anti_slave_0_readdata),    // SysID.readdata
		.avs_SysID_address     (basic_sysid_0_sysid_translator_avalon_anti_slave_0_address),     //      .address
		.avs_SysID_read        (basic_sysid_0_sysid_translator_avalon_anti_slave_0_read),        //      .read
		.avs_SysID_waitrequest (basic_sysid_0_sysid_translator_avalon_anti_slave_0_waitrequest)  //      .waitrequest
	);

	test_RegRW32 test_regrw32_0 (
		.rsi_MRST_reset       (qsys_serial_host_0_mrst_reset),                                  // MRST.reset
		.csi_MCLK_clk         (qsys_serial_host_0_mclk_clk),                                    // MCLK.clk
		.avs_test_writedata   (test_regrw32_0_test_translator_avalon_anti_slave_0_writedata),   // test.writedata
		.avs_test_readdata    (test_regrw32_0_test_translator_avalon_anti_slave_0_readdata),    //     .readdata
		.avs_test_byteenable  (test_regrw32_0_test_translator_avalon_anti_slave_0_byteenable),  //     .byteenable
		.avs_test_write       (test_regrw32_0_test_translator_avalon_anti_slave_0_write),       //     .write
		.avs_test_read        (test_regrw32_0_test_translator_avalon_anti_slave_0_read),        //     .read
		.avs_test_waitrequest (test_regrw32_0_test_translator_avalon_anti_slave_0_waitrequest)  //     .waitrequest
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (8),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (10),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (1),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (0),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) qsys_serial_host_0_m1_translator (
		.clk                   (qsys_serial_host_0_mclk_clk),                                              //                       clk.clk
		.reset                 (qsys_serial_host_0_mrst_reset),                                            //                     reset.reset
		.uav_address           (qsys_serial_host_0_m1_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (qsys_serial_host_0_m1_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (qsys_serial_host_0_m1_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (qsys_serial_host_0_m1_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (qsys_serial_host_0_m1_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (qsys_serial_host_0_m1_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (qsys_serial_host_0_m1_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (qsys_serial_host_0_m1_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (qsys_serial_host_0_m1_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (qsys_serial_host_0_m1_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (qsys_serial_host_0_m1_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (qsys_serial_host_0_m1_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (qsys_serial_host_0_m1_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (qsys_serial_host_0_m1_byteenable),                                         //                          .byteenable
		.av_begintransfer      (qsys_serial_host_0_m1_begintransfer),                                      //                          .begintransfer
		.av_read               (qsys_serial_host_0_m1_read),                                               //                          .read
		.av_readdata           (qsys_serial_host_0_m1_readdata),                                           //                          .readdata
		.av_readdatavalid      (qsys_serial_host_0_m1_readdatavalid),                                      //                          .readdatavalid
		.av_write              (qsys_serial_host_0_m1_write),                                              //                          .write
		.av_writedata          (qsys_serial_host_0_m1_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                     //               (terminated)
		.av_chipselect         (1'b0),                                                                     //               (terminated)
		.av_lock               (1'b0),                                                                     //               (terminated)
		.av_debugaccess        (1'b0),                                                                     //               (terminated)
		.uav_clken             (),                                                                         //               (terminated)
		.av_clken              (1'b1)                                                                      //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) basic_sysid_0_sysid_translator (
		.clk                   (qsys_serial_host_0_mclk_clk),                                                    //                      clk.clk
		.reset                 (qsys_serial_host_0_mrst_reset),                                                  //                    reset.reset
		.uav_address           (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (basic_sysid_0_sysid_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_read               (basic_sysid_0_sysid_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (basic_sysid_0_sysid_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (basic_sysid_0_sysid_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_write              (),                                                                               //              (terminated)
		.av_writedata          (),                                                                               //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_byteenable         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.av_chipselect         (),                                                                               //              (terminated)
		.av_clken              (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) test_regrw32_0_test_translator (
		.clk                   (qsys_serial_host_0_mclk_clk),                                                    //                      clk.clk
		.reset                 (qsys_serial_host_0_mrst_reset),                                                  //                    reset.reset
		.uav_address           (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (test_regrw32_0_test_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (test_regrw32_0_test_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (test_regrw32_0_test_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (test_regrw32_0_test_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (test_regrw32_0_test_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (test_regrw32_0_test_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                               //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.av_chipselect         (),                                                                               //              (terminated)
		.av_clken              (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (72),
		.PKT_PROTECTION_L          (70),
		.PKT_BEGIN_BURST           (65),
		.PKT_BURSTWRAP_H           (57),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BURST_SIZE_H          (60),
		.PKT_BURST_SIZE_L          (58),
		.PKT_BURST_TYPE_H          (62),
		.PKT_BURST_TYPE_L          (61),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_TRANS_EXCLUSIVE       (51),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (67),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (68),
		.PKT_DEST_ID_L             (68),
		.PKT_THREAD_ID_H           (69),
		.PKT_THREAD_ID_L           (69),
		.PKT_CACHE_H               (76),
		.PKT_CACHE_L               (73),
		.PKT_DATA_SIDEBAND_H       (64),
		.PKT_DATA_SIDEBAND_L       (64),
		.PKT_QOS_H                 (66),
		.PKT_QOS_L                 (66),
		.PKT_ADDR_SIDEBAND_H       (63),
		.PKT_ADDR_SIDEBAND_L       (63),
		.ST_DATA_W                 (79),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent (
		.clk              (qsys_serial_host_0_mclk_clk),                                                       //       clk.clk
		.reset            (qsys_serial_host_0_mrst_reset),                                                     // clk_reset.reset
		.av_address       (qsys_serial_host_0_m1_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (qsys_serial_host_0_m1_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (qsys_serial_host_0_m1_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (qsys_serial_host_0_m1_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (qsys_serial_host_0_m1_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (qsys_serial_host_0_m1_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (qsys_serial_host_0_m1_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (qsys_serial_host_0_m1_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (qsys_serial_host_0_m1_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (qsys_serial_host_0_m1_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (qsys_serial_host_0_m1_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                             //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                              //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                           //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                     //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                       //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                              //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (65),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (67),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (68),
		.PKT_DEST_ID_L             (68),
		.PKT_BURSTWRAP_H           (57),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (72),
		.PKT_PROTECTION_L          (70),
		.PKT_RESPONSE_STATUS_H     (78),
		.PKT_RESPONSE_STATUS_L     (77),
		.PKT_BURST_SIZE_H          (60),
		.PKT_BURST_SIZE_L          (58),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (79),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent (
		.clk                     (qsys_serial_host_0_mclk_clk),                                                              //             clk.clk
		.reset                   (qsys_serial_host_0_mrst_reset),                                                            //       clk_reset.reset
		.m0_address              (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src0_ready),                                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_src0_valid),                                                                //                .valid
		.cp_data                 (cmd_xbar_demux_src0_data),                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_src0_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src0_endofpacket),                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src0_channel),                                                              //                .channel
		.rf_sink_ready           (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (80),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (qsys_serial_host_0_mclk_clk),                                                              //       clk.clk
		.reset             (qsys_serial_host_0_mrst_reset),                                                            // clk_reset.reset
		.in_data           (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (65),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (67),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (68),
		.PKT_DEST_ID_L             (68),
		.PKT_BURSTWRAP_H           (57),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (72),
		.PKT_PROTECTION_L          (70),
		.PKT_RESPONSE_STATUS_H     (78),
		.PKT_RESPONSE_STATUS_L     (77),
		.PKT_BURST_SIZE_H          (60),
		.PKT_BURST_SIZE_L          (58),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (79),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) test_regrw32_0_test_translator_avalon_universal_slave_0_agent (
		.clk                     (qsys_serial_host_0_mclk_clk),                                                              //             clk.clk
		.reset                   (qsys_serial_host_0_mrst_reset),                                                            //       clk_reset.reset
		.m0_address              (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src1_ready),                                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_src1_valid),                                                                //                .valid
		.cp_data                 (cmd_xbar_demux_src1_data),                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_src1_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src1_endofpacket),                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src1_channel),                                                              //                .channel
		.rf_sink_ready           (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (80),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (qsys_serial_host_0_mclk_clk),                                                              //       clk.clk
		.reset             (qsys_serial_host_0_mrst_reset),                                                            // clk_reset.reset
		.in_data           (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	mse_addr_router addr_router (
		.sink_ready         (qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (qsys_serial_host_0_mclk_clk),                                                       //       clk.clk
		.reset              (qsys_serial_host_0_mrst_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_src_valid),                                                             //          .valid
		.src_data           (addr_router_src_data),                                                              //          .data
		.src_channel        (addr_router_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                        //          .endofpacket
	);

	mse_id_router id_router (
		.sink_ready         (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (basic_sysid_0_sysid_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (qsys_serial_host_0_mclk_clk),                                                    //       clk.clk
		.reset              (qsys_serial_host_0_mrst_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                            //       src.ready
		.src_valid          (id_router_src_valid),                                                            //          .valid
		.src_data           (id_router_src_data),                                                             //          .data
		.src_channel        (id_router_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                       //          .endofpacket
	);

	mse_id_router id_router_001 (
		.sink_ready         (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (test_regrw32_0_test_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (qsys_serial_host_0_mclk_clk),                                                    //       clk.clk
		.reset              (qsys_serial_host_0_mrst_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                        //       src.ready
		.src_valid          (id_router_001_src_valid),                                                        //          .valid
		.src_data           (id_router_001_src_data),                                                         //          .data
		.src_channel        (id_router_001_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                   //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (68),
		.PKT_DEST_ID_L             (68),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (79),
		.ST_CHANNEL_W              (2),
		.VALID_WIDTH               (2),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (qsys_serial_host_0_mclk_clk),    //       clk.clk
		.reset                  (qsys_serial_host_0_mrst_reset),  // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	mse_cmd_xbar_demux cmd_xbar_demux (
		.clk                (qsys_serial_host_0_mclk_clk),       //        clk.clk
		.reset              (qsys_serial_host_0_mrst_reset),     //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket)    //           .endofpacket
	);

	mse_rsp_xbar_demux rsp_xbar_demux (
		.clk                (qsys_serial_host_0_mclk_clk),       //       clk.clk
		.reset              (qsys_serial_host_0_mrst_reset),     // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)    //          .endofpacket
	);

	mse_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (qsys_serial_host_0_mclk_clk),           //       clk.clk
		.reset              (qsys_serial_host_0_mrst_reset),         // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	mse_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (qsys_serial_host_0_mclk_clk),           //       clk.clk
		.reset               (qsys_serial_host_0_mrst_reset),         // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

endmodule
