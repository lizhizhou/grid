// mse.v

// Generated using ACDS version 12.1sp1 243 at 2013.07.08.21:26:37

`timescale 1 ps / 1 ps
module mse (
		output wire  qsys_serial_host_0_sdo,   // qsys_serial_host_0.sdo
		input  wire  qsys_serial_host_0_sdi,   //                   .sdi
		input  wire  qsys_serial_host_0_clk,   //                   .clk
		input  wire  qsys_serial_host_0_sle,   //                   .sle
		output wire  qsys_serial_host_0_srdy,  //                   .srdy
		input  wire  qsys_serial_host_0_reset  //                   .reset
	);

	wire         qsys_serial_host_0_mrst_reset;                                            // qsys_serial_host_0:rso_MRST_reset -> [basic_SysID_0:rsi_MRST_reset, basic_SysID_0_SysID_translator:reset, qsys_serial_host_0_m1_translator:reset]
	wire         qsys_serial_host_0_mclk_clk;                                              // qsys_serial_host_0:cso_MCLK_clk -> [basic_SysID_0:csi_MCLK_clk, basic_SysID_0_SysID_translator:clk, qsys_serial_host_0_m1_translator:clk]
	wire         qsys_serial_host_0_m1_waitrequest;                                        // qsys_serial_host_0_m1_translator:av_waitrequest -> qsys_serial_host_0:avm_M1_waitrequest
	wire   [7:0] qsys_serial_host_0_m1_address;                                            // qsys_serial_host_0:avm_M1_address -> qsys_serial_host_0_m1_translator:av_address
	wire  [31:0] qsys_serial_host_0_m1_writedata;                                          // qsys_serial_host_0:avm_M1_writedata -> qsys_serial_host_0_m1_translator:av_writedata
	wire         qsys_serial_host_0_m1_write;                                              // qsys_serial_host_0:avm_M1_write -> qsys_serial_host_0_m1_translator:av_write
	wire         qsys_serial_host_0_m1_read;                                               // qsys_serial_host_0:avm_M1_read -> qsys_serial_host_0_m1_translator:av_read
	wire  [31:0] qsys_serial_host_0_m1_readdata;                                           // qsys_serial_host_0_m1_translator:av_readdata -> qsys_serial_host_0:avm_M1_readdata
	wire         qsys_serial_host_0_m1_begintransfer;                                      // qsys_serial_host_0:avm_M1_begintransfer -> qsys_serial_host_0_m1_translator:av_begintransfer
	wire         qsys_serial_host_0_m1_readdatavalid;                                      // qsys_serial_host_0_m1_translator:av_readdatavalid -> qsys_serial_host_0:avm_M1_readdatavalid
	wire   [3:0] qsys_serial_host_0_m1_byteenable;                                         // qsys_serial_host_0:avm_M1_byteenable -> qsys_serial_host_0_m1_translator:av_byteenable
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_waitrequest;   // basic_SysID_0_SysID_translator:uav_waitrequest -> qsys_serial_host_0_m1_translator:uav_waitrequest
	wire   [2:0] qsys_serial_host_0_m1_translator_avalon_universal_master_0_burstcount;    // qsys_serial_host_0_m1_translator:uav_burstcount -> basic_SysID_0_SysID_translator:uav_burstcount
	wire  [31:0] qsys_serial_host_0_m1_translator_avalon_universal_master_0_writedata;     // qsys_serial_host_0_m1_translator:uav_writedata -> basic_SysID_0_SysID_translator:uav_writedata
	wire   [9:0] qsys_serial_host_0_m1_translator_avalon_universal_master_0_address;       // qsys_serial_host_0_m1_translator:uav_address -> basic_SysID_0_SysID_translator:uav_address
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_lock;          // qsys_serial_host_0_m1_translator:uav_lock -> basic_SysID_0_SysID_translator:uav_lock
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_write;         // qsys_serial_host_0_m1_translator:uav_write -> basic_SysID_0_SysID_translator:uav_write
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_read;          // qsys_serial_host_0_m1_translator:uav_read -> basic_SysID_0_SysID_translator:uav_read
	wire  [31:0] qsys_serial_host_0_m1_translator_avalon_universal_master_0_readdata;      // basic_SysID_0_SysID_translator:uav_readdata -> qsys_serial_host_0_m1_translator:uav_readdata
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_debugaccess;   // qsys_serial_host_0_m1_translator:uav_debugaccess -> basic_SysID_0_SysID_translator:uav_debugaccess
	wire   [3:0] qsys_serial_host_0_m1_translator_avalon_universal_master_0_byteenable;    // qsys_serial_host_0_m1_translator:uav_byteenable -> basic_SysID_0_SysID_translator:uav_byteenable
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_readdatavalid; // basic_SysID_0_SysID_translator:uav_readdatavalid -> qsys_serial_host_0_m1_translator:uav_readdatavalid
	wire         basic_sysid_0_sysid_translator_avalon_anti_slave_0_waitrequest;           // basic_SysID_0:avs_SysID_waitrequest -> basic_SysID_0_SysID_translator:av_waitrequest
	wire   [1:0] basic_sysid_0_sysid_translator_avalon_anti_slave_0_address;               // basic_SysID_0_SysID_translator:av_address -> basic_SysID_0:avs_SysID_address
	wire         basic_sysid_0_sysid_translator_avalon_anti_slave_0_read;                  // basic_SysID_0_SysID_translator:av_read -> basic_SysID_0:avs_SysID_read
	wire  [31:0] basic_sysid_0_sysid_translator_avalon_anti_slave_0_readdata;              // basic_SysID_0:avs_SysID_readdata -> basic_SysID_0_SysID_translator:av_readdata

	qsys_serial_host #(
		.initial_state (9'b000000000)
	) qsys_serial_host_0 (
		.rso_MRST_reset       (qsys_serial_host_0_mrst_reset),       //        mrst.reset
		.cso_MCLK_clk         (qsys_serial_host_0_mclk_clk),         //        mclk.clk
		.avm_M1_writedata     (qsys_serial_host_0_m1_writedata),     //          m1.writedata
		.avm_M1_readdata      (qsys_serial_host_0_m1_readdata),      //            .readdata
		.avm_M1_address       (qsys_serial_host_0_m1_address),       //            .address
		.avm_M1_byteenable    (qsys_serial_host_0_m1_byteenable),    //            .byteenable
		.avm_M1_write         (qsys_serial_host_0_m1_write),         //            .write
		.avm_M1_read          (qsys_serial_host_0_m1_read),          //            .read
		.avm_M1_begintransfer (qsys_serial_host_0_m1_begintransfer), //            .begintransfer
		.avm_M1_readdatavalid (qsys_serial_host_0_m1_readdatavalid), //            .readdatavalid
		.avm_M1_waitrequest   (qsys_serial_host_0_m1_waitrequest),   //            .waitrequest
		.sdo                  (qsys_serial_host_0_sdo),              // conduit_end.export
		.sdi                  (qsys_serial_host_0_sdi),              //            .export
		.clk                  (qsys_serial_host_0_clk),              //            .export
		.sle                  (qsys_serial_host_0_sle),              //            .export
		.srdy                 (qsys_serial_host_0_srdy),             //            .export
		.reset                (qsys_serial_host_0_reset)             //            .export
	);

	basic_SysID basic_sysid_0 (
		.rsi_MRST_reset        (qsys_serial_host_0_mrst_reset),                                  //  MRST.reset
		.csi_MCLK_clk          (qsys_serial_host_0_mclk_clk),                                    //  MCLK.clk
		.avs_SysID_readdata    (basic_sysid_0_sysid_translator_avalon_anti_slave_0_readdata),    // SysID.readdata
		.avs_SysID_address     (basic_sysid_0_sysid_translator_avalon_anti_slave_0_address),     //      .address
		.avs_SysID_read        (basic_sysid_0_sysid_translator_avalon_anti_slave_0_read),        //      .read
		.avs_SysID_waitrequest (basic_sysid_0_sysid_translator_avalon_anti_slave_0_waitrequest)  //      .waitrequest
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (8),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (10),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (1),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (0),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) qsys_serial_host_0_m1_translator (
		.clk                   (qsys_serial_host_0_mclk_clk),                                              //                       clk.clk
		.reset                 (qsys_serial_host_0_mrst_reset),                                            //                     reset.reset
		.uav_address           (qsys_serial_host_0_m1_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (qsys_serial_host_0_m1_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (qsys_serial_host_0_m1_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (qsys_serial_host_0_m1_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (qsys_serial_host_0_m1_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (qsys_serial_host_0_m1_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (qsys_serial_host_0_m1_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (qsys_serial_host_0_m1_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (qsys_serial_host_0_m1_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (qsys_serial_host_0_m1_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (qsys_serial_host_0_m1_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (qsys_serial_host_0_m1_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (qsys_serial_host_0_m1_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (qsys_serial_host_0_m1_byteenable),                                         //                          .byteenable
		.av_begintransfer      (qsys_serial_host_0_m1_begintransfer),                                      //                          .begintransfer
		.av_read               (qsys_serial_host_0_m1_read),                                               //                          .read
		.av_readdata           (qsys_serial_host_0_m1_readdata),                                           //                          .readdata
		.av_readdatavalid      (qsys_serial_host_0_m1_readdatavalid),                                      //                          .readdatavalid
		.av_write              (qsys_serial_host_0_m1_write),                                              //                          .write
		.av_writedata          (qsys_serial_host_0_m1_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                     //               (terminated)
		.av_chipselect         (1'b0),                                                                     //               (terminated)
		.av_lock               (1'b0),                                                                     //               (terminated)
		.av_debugaccess        (1'b0),                                                                     //               (terminated)
		.uav_clken             (),                                                                         //               (terminated)
		.av_clken              (1'b1)                                                                      //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) basic_sysid_0_sysid_translator (
		.clk                   (qsys_serial_host_0_mclk_clk),                                              //                      clk.clk
		.reset                 (qsys_serial_host_0_mrst_reset),                                            //                    reset.reset
		.uav_address           (qsys_serial_host_0_m1_translator_avalon_universal_master_0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (qsys_serial_host_0_m1_translator_avalon_universal_master_0_burstcount),    //                         .burstcount
		.uav_read              (qsys_serial_host_0_m1_translator_avalon_universal_master_0_read),          //                         .read
		.uav_write             (qsys_serial_host_0_m1_translator_avalon_universal_master_0_write),         //                         .write
		.uav_waitrequest       (qsys_serial_host_0_m1_translator_avalon_universal_master_0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (qsys_serial_host_0_m1_translator_avalon_universal_master_0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (qsys_serial_host_0_m1_translator_avalon_universal_master_0_byteenable),    //                         .byteenable
		.uav_readdata          (qsys_serial_host_0_m1_translator_avalon_universal_master_0_readdata),      //                         .readdata
		.uav_writedata         (qsys_serial_host_0_m1_translator_avalon_universal_master_0_writedata),     //                         .writedata
		.uav_lock              (qsys_serial_host_0_m1_translator_avalon_universal_master_0_lock),          //                         .lock
		.uav_debugaccess       (qsys_serial_host_0_m1_translator_avalon_universal_master_0_debugaccess),   //                         .debugaccess
		.av_address            (basic_sysid_0_sysid_translator_avalon_anti_slave_0_address),               //      avalon_anti_slave_0.address
		.av_read               (basic_sysid_0_sysid_translator_avalon_anti_slave_0_read),                  //                         .read
		.av_readdata           (basic_sysid_0_sysid_translator_avalon_anti_slave_0_readdata),              //                         .readdata
		.av_waitrequest        (basic_sysid_0_sysid_translator_avalon_anti_slave_0_waitrequest),           //                         .waitrequest
		.av_write              (),                                                                         //              (terminated)
		.av_writedata          (),                                                                         //              (terminated)
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

endmodule
