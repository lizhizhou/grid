library verilog;
use verilog.vl_types.all;
entity port_io_interface_sim is
end port_io_interface_sim;
